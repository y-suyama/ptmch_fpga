//==================================================================================================
//  Company name        : 
//  Date                : 
//  File Name           : max10_10m08_top.v
//  Project Name        : 
//  Coding              : suyama
//  Rev.                : 1.0
//
//==================================================================================================
// Import
//==================================================================================================
// None
//==================================================================================================
// Module
//==================================================================================================
module max10_10m08_top(
    // Clock, Reset
    input  logic         CLK50M,
    input  logic         RESET_N,
    // SPI Signal
    input  logic         SPI_CS,
    input  logic         SPI_CLK,
    input  logic         SPI_MOSI,
    output logic [ 3: 0] TRG_PLS
);
//=================================================================
//  Internal Signal
//=================================================================
    logic  w_clk160m;
//=================================================================
//  output Port
//=================================================================
//==================================================================================================
//  Structural coding
//==================================================================================================

nios2_system u0(
    .clock_clk                    (CLK50M),
    .reset_n_reset_n              (RESET_N),
    .altpll_0_c1_clk              (w_clk160m)
   );

ptmch_top ptmch_inst(
    // Reset/Clock
    .RESET_N(RESET_N),
    .CLK160M(w_clk160m),
    // SPI Interface
    .SPI_CS(SPI_CS),
    .SPI_CLK(SPI_CLK),
    .SPI_MOSI(SPI_MOSI),
    .TRG_PLS(TRG_PLS)
);

endmodule
