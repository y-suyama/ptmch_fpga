//==================================================================================================
//  Company name        : 
//  Date                : 
//  File Name           : ptmch_top.sv
//  Project Name        : 
//  Coding              : suyama
//  Rev.                : 1.0
//
//==================================================================================================
// Import
//==================================================================================================
// None
//==================================================================================================
// Module
//==================================================================================================
module ptmch_top(
    // Reset/Clock
    input  logic        RESET_N,
    input  logic        CLK200M,
 //   input  logic        CLK100M,
    // SPI Interface
    input  logic        SPI_CS,
    input  logic        SPI_CLK,
    input  logic        SPI_MOSI,
    output logic        TRG_PLS
);
//==================================================================================================
//  PARAMETER declarations
//==================================================================================================
//    parameter p_addrexpander   = 16'h3000;
//==================================================================================================
//  Internal Signal
//==================================================================================================

//==================================================================================================
//  output Port
//==================================================================================================

//==================================================================================================
//  Structural coding
//==================================================================================================

ptmch_trg trg_inst(
    .RESET_N(RESET_N),
    .CLK200M(CLK200M),
    .SPI_CS(SPI_CS),
    .SPI_CLK(SPI_CLK),
    .SPI_MOSI(SPI_MOSI),
    .TRG_PLS(TRG_PLS)
);

endmodule
