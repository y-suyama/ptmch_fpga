
module nios2_system (
	altpll_0_c1_clk,
	clock_clk,
	reset_n_reset_n);	

	output		altpll_0_c1_clk;
	input		clock_clk;
	input		reset_n_reset_n;
endmodule
